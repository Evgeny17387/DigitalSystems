module alu64bit_test;







endmodule
